`include "define.v"

module fake_mem_if(
    input wire reset,

    input wire [`MemAddrBus] pc,
    output reg [`InstBus] inst
);

    always @(*) begin
        if (reset == 1) begin
            inst <= 0;
        end else begin
            case (pc)
                0: inst <= 32'b0000000_11011_10110_011_01011_0110011;
                4: inst <= 32'b0000000_11101_11011_100_11001_0110011;
                8: inst <= 32'b100111011001_00101_010_10010_0010011;
                12: inst <= 32'b011110000110_10001_000_10010_0010011;
                16: inst <= 32'b0000000_10101_11000_100_01100_0110011;
                20: inst <= 32'b0000000_00111_11000_011_10000_0110011;
                24: inst <= 32'b0000000_00000_00101_101_01000_0110011;
                28: inst <= 32'b001101000001_11000_000_10010_0010011;
                32: inst <= 32'b110100000100_11100_011_10101_0010011;
                36: inst <= 32'b0000000_00111_01001_101_00110_0110011;
                40: inst <= 32'b0000000_11000_11101_001_10010_0010011;
                44: inst <= 32'b011011100110_11010_011_11000_0010011;
                48: inst <= 32'b0100000_11000_00101_101_10010_0010011;
                52: inst <= 32'b0000000_00010_10001_111_10100_0110011;
                56: inst <= 32'b110000010010_10111_100_11100_0010011;
                60: inst <= 32'b0100000_00101_11100_000_10000_0110011;
                64: inst <= 32'b101110101101_11111_100_01101_0010011;
                68: inst <= 32'b0000000_11000_01111_110_00001_0110011;
                72: inst <= 32'b0000000_00000_00011_110_01011_0110011;
                76: inst <= 32'b0000000_11011_01001_101_01111_0010011;
                80: inst <= 32'b0000000_01111_00101_101_10011_0010011;
                84: inst <= 32'b0100000_11100_01101_101_11100_0010011;
                88: inst <= 32'b0000000_01010_01001_110_11100_0110011;
                92: inst <= 32'b0000000_10101_00101_111_10011_0110011;
                96: inst <= 32'b011101111010_00110_110_11000_0010011;
                100: inst <= 32'b0100000_01011_01011_101_01110_0110011;
                104: inst <= 32'b0000000_01001_10011_101_01011_0110011;
                108: inst <= 32'b101000111100_10000_011_10010_0010011;
                112: inst <= 32'b0000000_10110_11111_001_10010_0110011;
                116: inst <= 32'b0000000_00110_10000_100_11101_0110011;
                120: inst <= 32'b0000000_00111_10010_101_01011_0010011;
                124: inst <= 32'b000101100110_10001_110_11011_0010011;
                128: inst <= 32'b100001111010_00011_110_11001_0010011;
                132: inst <= 32'b0000000_00011_00000_001_11000_0110011;
                136: inst <= 32'b001101010110_01010_010_00011_0010011;
                140: inst <= 32'b0000000_01110_01011_101_11101_0110011;
                144: inst <= 32'b0000000_00011_00111_110_10011_0110011;
                148: inst <= 32'b0000000_10110_00100_010_01101_0110011;
                152: inst <= 32'b110101011011_01111_110_10101_0010011;
                156: inst <= 32'b0000000_00100_11100_011_00101_0110011;
                160: inst <= 32'b0000000_11110_11010_001_01110_0010011;
                164: inst <= 32'b0000000_00011_01110_101_01010_0110011;
                168: inst <= 32'b0000000_11000_11101_010_10011_0110011;
                172: inst <= 32'b111110111110_10011_010_11000_0010011;
                176: inst <= 32'b001001001000_11001_100_11001_0010011;
                180: inst <= 32'b0000000_01100_01000_101_10101_0010011;
                184: inst <= 32'b0000000_10101_10101_000_00001_0110011;
                188: inst <= 32'b010011101111_10101_111_00110_0010011;
                192: inst <= 32'b0000000_11101_01011_100_11011_0110011;
                196: inst <= 32'b001111001000_01101_011_11100_0010011;
                200: inst <= 32'b100100101110_11110_100_10100_0010011;
                204: inst <= 32'b0100000_01110_01101_101_01111_0010011;
                208: inst <= 32'b0000000_01100_00011_011_00001_0110011;
                212: inst <= 32'b0100000_01011_01101_000_10101_0110011;
                216: inst <= 32'b101101010111_11110_111_01000_0010011;
                220: inst <= 32'b0000000_01111_00001_001_11011_0110011;
                224: inst <= 32'b011001111001_01111_000_11110_0010011;
                228: inst <= 32'b011000110111_10010_010_10010_0010011;
                232: inst <= 32'b0000000_10000_01010_010_00100_0110011;
                236: inst <= 32'b0100000_10011_01000_101_10011_0010011;
                240: inst <= 32'b101111010011_00001_011_00110_0010011;
                244: inst <= 32'b0100000_11100_01001_101_10110_0110011;
                248: inst <= 32'b0100000_11000_00000_101_00001_0110011;
                252: inst <= 32'b0000000_01011_01100_011_00110_0110011;
                256: inst <= 32'b011101000101_11001_100_11101_0010011;
                260: inst <= 32'b010100111111_01010_110_01011_0010011;
                264: inst <= 32'b110111001011_10111_010_00101_0010011;
                268: inst <= 32'b010101011101_01100_100_00110_0010011;
                272: inst <= 32'b0100000_01001_01100_000_01010_0110011;
                276: inst <= 32'b010010001010_01100_000_11100_0010011;
                280: inst <= 32'b0000000_11110_11000_010_01101_0110011;
                284: inst <= 32'b0000000_11011_01110_001_00100_0110011;
                288: inst <= 32'b0000000_10010_00111_011_00111_0110011;
                292: inst <= 32'b0100000_10000_01100_101_00101_0110011;
                296: inst <= 32'b0100000_00010_11100_000_01111_0110011;
                300: inst <= 32'b0000000_00010_00001_100_00110_0110011;
                304: inst <= 32'b000100000010_11111_010_01101_0010011;
                308: inst <= 32'b011110011111_00111_010_11001_0010011;
                312: inst <= 32'b0000000_01011_00010_010_01010_0110011;
                316: inst <= 32'b110110101111_10011_111_10010_0010011;
                320: inst <= 32'b0000000_00101_00111_010_01001_0110011;
                324: inst <= 32'b011110110111_10100_000_01111_0010011;
                328: inst <= 32'b0000000_10010_10000_111_00001_0110011;
                332: inst <= 32'b0000000_01001_00010_101_00001_0010011;
                336: inst <= 32'b101101001010_11001_100_10101_0010011;
                340: inst <= 32'b0000000_10111_11101_001_11110_0110011;
                344: inst <= 32'b0000000_01100_00011_001_10001_0010011;
                348: inst <= 32'b0000000_00110_00010_010_11001_0110011;
                352: inst <= 32'b0000000_00011_10011_010_10101_0110011;
                356: inst <= 32'b0000000_11111_00011_001_01111_0110011;
                360: inst <= 32'b0000000_10000_11110_100_10100_0110011;
                364: inst <= 32'b101111101000_01111_110_11101_0010011;
                368: inst <= 32'b111111000111_00110_111_11011_0010011;
                372: inst <= 32'b0000000_11111_01011_111_01001_0110011;
                376: inst <= 32'b100000101100_10011_011_11110_0010011;
                380: inst <= 32'b011010011000_00010_110_11110_0010011;
                384: inst <= 32'b001101001001_00101_011_01010_0010011;
                388: inst <= 32'b0000000_11001_11111_101_01010_0010011;
                392: inst <= 32'b0000000_00010_10000_011_11011_0110011;
                396: inst <= 32'b0100000_01111_11001_101_10011_0110011;
                400: inst <= 32'b110111111000_00011_111_01011_0010011;
                404: inst <= 32'b0000000_11110_01000_101_01000_0010011;
                408: inst <= 32'b001001101001_01001_000_00100_0010011;
                412: inst <= 32'b0000000_11100_00011_001_10000_0010011;
                416: inst <= 32'b011110100110_11100_111_11001_0010011;
                420: inst <= 32'b0000000_10011_00101_001_00110_0110011;
                424: inst <= 32'b0000000_10100_11010_110_00110_0110011;
                428: inst <= 32'b0000000_11101_01111_001_11011_0010011;
                432: inst <= 32'b0000000_01101_00111_011_10000_0110011;
                436: inst <= 32'b0100000_00111_10001_101_11101_0010011;
                440: inst <= 32'b0000000_00001_10100_100_11100_0110011;
                444: inst <= 32'b0000000_10100_11000_101_10001_0010011;
                448: inst <= 32'b0100000_11010_11010_101_01111_0010011;
                452: inst <= 32'b0000000_10100_01001_010_10001_0110011;
                456: inst <= 32'b0000000_01010_11111_111_00101_0110011;
                460: inst <= 32'b0000000_11011_10110_001_10011_0010011;
                464: inst <= 32'b0000000_10000_10100_100_01101_0110011;
                468: inst <= 32'b0100000_00110_00011_101_00110_0110011;
                472: inst <= 32'b0100000_11101_10100_101_10011_0110011;
                476: inst <= 32'b0000000_10100_10011_101_10101_0110011;
                480: inst <= 32'b0100000_00001_01101_000_10000_0110011;
                484: inst <= 32'b0100000_11010_01101_101_10011_0010011;
                488: inst <= 32'b100100111000_10111_111_10001_0010011;
                492: inst <= 32'b110100010111_11011_000_01011_0010011;
                496: inst <= 32'b0100000_01001_01111_101_01100_0110011;
                500: inst <= 32'b0000000_00001_11100_101_00111_0110011;
                504: inst <= 32'b0000000_10001_11100_100_01101_0110011;
                508: inst <= 32'b0000000_11110_01010_101_00100_0010011;
                512: inst <= 32'b0000000_01110_10110_101_10001_0010011;
                516: inst <= 32'b0100000_10101_10010_000_00101_0110011;
                520: inst <= 32'b001111000011_10110_111_00110_0010011;
                524: inst <= 32'b0000000_11111_01100_100_11001_0110011;
                528: inst <= 32'b0000000_00001_10110_101_11101_0110011;
                532: inst <= 32'b111000100110_10001_110_10001_0010011;
                536: inst <= 32'b0000000_00001_01110_011_01100_0110011;
                540: inst <= 32'b0000000_01000_10011_111_01101_0110011;
                544: inst <= 32'b0000000_10110_01010_011_01010_0110011;
                548: inst <= 32'b101101001000_00010_110_11001_0010011;
                552: inst <= 32'b0000000_00111_00010_000_10100_0110011;
                556: inst <= 32'b0000000_01101_11100_110_10110_0110011;
                560: inst <= 32'b0000000_11000_10011_000_10000_0110011;
                564: inst <= 32'b0000000_00001_10100_110_00011_0110011;
                568: inst <= 32'b111100100100_11110_100_00111_0010011;
                572: inst <= 32'b0100000_01111_01101_101_10010_0010011;
                576: inst <= 32'b100000111011_11000_010_10000_0010011;
                580: inst <= 32'b0000000_11100_10101_101_01101_0110011;
                584: inst <= 32'b0000000_10000_11010_010_11100_0110011;
                588: inst <= 32'b0000000_00101_01001_100_01111_0110011;
                592: inst <= 32'b0000000_00001_00001_100_01011_0110011;
                596: inst <= 32'b0000000_11111_00100_001_10111_0110011;
                600: inst <= 32'b011001111011_10000_111_11111_0010011;
                604: inst <= 32'b0000000_11010_10010_001_10010_0110011;
                608: inst <= 32'b0000000_01010_11010_111_01111_0110011;
                612: inst <= 32'b0000000_00011_11101_011_10000_0110011;
                616: inst <= 32'b0000000_01010_00100_001_01000_0010011;
                620: inst <= 32'b0000000_10101_10000_100_01000_0110011;
                624: inst <= 32'b100010000101_00011_110_01110_0010011;
                628: inst <= 32'b010010000100_10111_000_11111_0010011;
                632: inst <= 32'b0100000_01101_00011_000_11010_0110011;
                636: inst <= 32'b000111100101_10001_000_10010_0010011;
                640: inst <= 32'b100101000101_00110_110_10001_0010011;
                644: inst <= 32'b0000000_11110_00010_011_01101_0110011;
                648: inst <= 32'b0100000_11010_10111_101_10101_0110011;
                652: inst <= 32'b0000000_00011_00001_100_10110_0110011;
                656: inst <= 32'b0000000_01010_10001_100_10000_0110011;
                660: inst <= 32'b0000000_11010_10001_101_01111_0110011;
                664: inst <= 32'b011101100001_00111_111_11001_0010011;
                668: inst <= 32'b0000000_11100_10101_001_10001_0110011;
                672: inst <= 32'b110110101101_00111_010_11100_0010011;
                676: inst <= 32'b0000000_10110_11110_001_10110_0010011;
                680: inst <= 32'b0000000_01101_10000_100_11111_0110011;
                684: inst <= 32'b010111100010_10111_000_01110_0010011;
                688: inst <= 32'b0000000_11111_01100_010_11111_0110011;
                692: inst <= 32'b0000000_00110_01111_011_01000_0110011;
                696: inst <= 32'b0000000_00001_01101_000_00110_0110011;
                700: inst <= 32'b011000101101_00010_100_11010_0010011;
                704: inst <= 32'b0100000_01111_00000_101_00101_0010011;
                708: inst <= 32'b0000000_00101_00011_001_11100_0010011;
                712: inst <= 32'b011010001111_11100_000_01001_0010011;
                716: inst <= 32'b111111001011_01001_000_01010_0010011;
                720: inst <= 32'b0000000_11001_01011_110_11100_0110011;
                724: inst <= 32'b0000000_00101_11110_011_10100_0110011;
                728: inst <= 32'b0100000_10001_11101_101_00010_0110011;
                732: inst <= 32'b0000000_01011_01110_010_10011_0110011;
                736: inst <= 32'b0000000_00111_00110_111_00111_0110011;
                740: inst <= 32'b001011100010_01001_011_01001_0010011;
                744: inst <= 32'b0100000_00000_11010_101_10100_0110011;
                748: inst <= 32'b0000000_00000_11110_111_01011_0110011;
                752: inst <= 32'b010100000110_00011_011_01110_0010011;
                756: inst <= 32'b0100000_00001_11101_101_10000_0010011;
                760: inst <= 32'b0100000_01100_10101_000_11111_0110011;
                764: inst <= 32'b0000000_00100_01010_101_11100_0010011;
                768: inst <= 32'b0000000_01111_01000_001_00101_0110011;
                772: inst <= 32'b0000000_01011_11000_001_10101_0010011;
                776: inst <= 32'b0100000_11000_11100_000_01001_0110011;
                780: inst <= 32'b100100111010_11100_110_01011_0010011;
                784: inst <= 32'b0000000_10000_00111_010_10011_0110011;
                788: inst <= 32'b101110101000_01101_010_10011_0010011;
                792: inst <= 32'b0000000_10010_01111_011_11000_0110011;
                796: inst <= 32'b0000000_00000_11000_110_11000_0110011;
                800: inst <= 32'b100100011011_10010_000_10111_0010011;
                804: inst <= 32'b011111011110_11110_000_01101_0010011;
                808: inst <= 32'b0100000_01101_10101_101_00100_0110011;
                812: inst <= 32'b0100000_00101_11100_000_10011_0110011;
                816: inst <= 32'b0000000_11100_00011_100_00010_0110011;
                820: inst <= 32'b0000000_10011_11100_100_11010_0110011;
                824: inst <= 32'b0100000_00110_00001_000_11011_0110011;
                828: inst <= 32'b0000000_01101_01100_110_11001_0110011;
                832: inst <= 32'b0000000_11000_01101_010_01110_0110011;
                836: inst <= 32'b0000000_00101_01010_101_01100_0010011;
                840: inst <= 32'b000001010011_10001_111_00011_0010011;
                844: inst <= 32'b0000000_00000_01000_100_00001_0110011;
                848: inst <= 32'b0000000_10110_11111_100_01010_0110011;
                852: inst <= 32'b001101000101_00000_111_10101_0010011;
                856: inst <= 32'b0000000_11000_10100_101_10011_0110011;
                860: inst <= 32'b0100000_10110_00011_101_11010_0010011;
                864: inst <= 32'b0000000_00010_10101_001_11000_0110011;
                868: inst <= 32'b0000000_11011_10110_111_00011_0110011;
                872: inst <= 32'b0000000_01001_00001_110_10111_0110011;
                876: inst <= 32'b0000000_00101_11100_011_01101_0110011;
                880: inst <= 32'b0000000_00111_01110_111_11010_0110011;
                884: inst <= 32'b0100000_00000_11000_000_00010_0110011;
                888: inst <= 32'b0000000_01110_11010_110_10101_0110011;
                892: inst <= 32'b0000000_00111_00010_010_11101_0110011;
                896: inst <= 32'b010010100110_01010_010_01000_0010011;
                900: inst <= 32'b0100000_00011_00011_101_00110_0110011;
                904: inst <= 32'b0000000_01010_11110_110_10111_0110011;
                908: inst <= 32'b0100000_11111_10111_101_10010_0110011;
                912: inst <= 32'b0000000_10111_00011_101_01111_0110011;
                916: inst <= 32'b0000000_11100_01010_111_00111_0110011;
                920: inst <= 32'b001010110011_00011_100_01101_0010011;
                924: inst <= 32'b100011001110_01010_100_01111_0010011;
                928: inst <= 32'b0000000_00001_11000_001_11010_0010011;
                932: inst <= 32'b0000000_01000_11100_101_11100_0010011;
                936: inst <= 32'b100110001011_01000_110_00011_0010011;
                940: inst <= 32'b100101001101_11010_110_01111_0010011;
                944: inst <= 32'b101100000100_10000_111_00001_0010011;
                948: inst <= 32'b0000000_10111_00000_101_01111_0010011;
                952: inst <= 32'b0000000_10010_01101_111_11010_0110011;
                956: inst <= 32'b0000000_10011_10100_101_11000_0010011;
                960: inst <= 32'b0000000_00010_11000_001_01001_0110011;
                964: inst <= 32'b001101001101_10101_110_01110_0010011;
                968: inst <= 32'b010000111010_10010_100_01011_0010011;
                972: inst <= 32'b011110011011_01000_111_00001_0010011;
                976: inst <= 32'b0000000_11110_00001_010_01100_0110011;
                980: inst <= 32'b011111110010_01111_110_11000_0010011;
                984: inst <= 32'b100001110001_01010_111_00110_0010011;
                988: inst <= 32'b100011100110_01000_110_10000_0010011;
                992: inst <= 32'b010101100001_00000_011_01101_0010011;
                996: inst <= 32'b101001001100_10100_000_11001_0010011;
                default : inst <= 0;
            endcase
        end
    end

endmodule
